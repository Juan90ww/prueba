`timescale 1ns/1ps

module tb_top_divisor_debug;

    logic clk = 0;
    logic rst = 0;

    logic [3:0] fil = 4'hF;

    wire [3:0] col;
    wire [3:0] anodo;
    wire [6:0] seven;

    wire [7:0] A_debug;
    wire [7:0] B_debug;
    wire [6:0] Q_debug;
    wire [6:0] R_debug;
    wire       done_debug;

    // Clock 50 MHz
    always #10 clk = ~clk;

    // Instancia del módulo top
    top_divisor_debug dut (
        .clk(clk),
        .rst(rst),
        .fil(fil),
        .col(col),
        .anodo(anodo),
        .seven(seven),
        .A_bin_debug(A_debug),
        .B_bin_debug(B_debug),
        .Q_debug(Q_debug),
        .R_debug(R_debug),
        .div_done_debug(done_debug)
    );

    // =====================================================
    // ENVÍO DE NIBBLES (estable y robusto)
    // =====================================================
    task send_nibble(input [3:0] val);
        begin
            fil = 4'hF;
            repeat (5) @(posedge clk);

            fil = val;         // mandar nibble
            repeat (5) @(posedge clk);

            fil = 4'hF;        // volver a idle
            repeat (5) @(posedge clk);
        end
    endtask

    task send_hex(input [7:0] val);
        begin
            send_nibble(val[7:4]);   // nibble alto
            send_nibble(val[3:0]);   // nibble bajo
        end
    endtask

    // =====================================================
    // TEST
    // =====================================================
    initial begin
        $dumpfile("tb_top_divisor_debug.vcd");
        $dumpvars(0, tb_top_divisor_debug);

        // Reset inicial
        rst = 0;
        repeat(10) @(posedge clk);
        rst = 1;
        repeat(10) @(posedge clk);

        $display("\n=== TEST: A=0x45, B=0x07 ===");

        send_hex(8'h45);   // A = 69 decimal
        send_hex(8'h07);   // B = 7 decimal

        @(posedge done_debug);

        $display("A=%0d  B=%0d  Q=%0d  R=%0d",
                 A_debug, B_debug, Q_debug, R_debug);

        repeat(20) @(posedge clk);

        $display("\nFIN SIMULACIÓN");
        $finish;
    end

endmodule

